//============================================================================
// Copyright(c) 2022 , Inchi Technology Inc, All right reserved
// Company           : Inchi Technology .Inc
//============================================================================
// Project           :vpu
// File Name         :instr_if.sv
// Author            :=huangxiaogang
// Email             :=huangxiaogang@inchitech.com
// Called by         :
// Reversion History :2023-09-04 14:45:34
// Reversion:        1.0
//============================================================================
// Description       :
//============================================================================

`ifndef _INSTR_IF_SV_
`define _INSTR_IF_SV_

interface instr_if(input clk, input rst_n);

  // You could add properties and assertions, for example
  // property name 
  // ...
  // endproperty : name
  // label: assert property(name)

endinterface : instr_if

`endif // INSTR_IF_SV
